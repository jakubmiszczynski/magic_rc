Inverter Simulation
* this file edited to remove everything not in tt lib
.lib "/home/kuba/.volare/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

* instantiate the inverter
X1R ONE TWO VGND X1

.subckt X1 one two VSUBS

* NGSPICE file created from magic_rc.ext - technology: sky130A

*.subckt magic_rc
X0 TWO TWO VSUBS sky130_fd_pr__res_xhigh_po w=2e+06u l=3.5e+06u
X1 TWO ONE VSUBS sky130_fd_pr__res_xhigh_po w=4e+06u l=5e+06u
X2 ONE ONE VSUBS sky130_fd_pr__res_xhigh_po w=2e+06u l=3.5e+06u
C0 ONE TWO 0.05fF
C1 TWO VSUBS 0.59fF
C2 down VSUBS 0.07fF $ **FLOATING
C3 ONE VSUBS 0.63fF
.ends

*.ends

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

R TWO VGND 10000

* create pulse
Vin ONE VGND pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10p 2n 0

.control
run
set color0 = white
set color1 = black
plot ONE TWO
.endc

.end

