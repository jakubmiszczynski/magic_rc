.ends

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

R TWO VGND 10000

* create pulse
Vin ONE VGND pulse(0 1.8 1p 10p 10p 1n 2n)
.tran 10p 2n 0

.control
run
set color0 = white
set color1 = black
plot ONE TWO
.endc

.end

